module concatenate(
  
);

endmodule