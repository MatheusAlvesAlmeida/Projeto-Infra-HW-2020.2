module det_size (
  input  wire [1:0] DetSizeCtrl,
  input  wire [31:0] data_in,
  output wire [31:0] data_out,
);

  assign data_out = 

endmodule