module set_size (
  input  wire [1:0] SetSizeCtrl,
  output wire [27:0] data_out,
);

  assign data_out = 

endmodule