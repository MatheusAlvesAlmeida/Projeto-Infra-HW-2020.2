module divisor(
    input wire clock,
    input wire reset,
    input wire multOrDiv,
    input signed [31:0] A,
    input signed [31:0] B,
    output reg [31:0] hi, 
    output reg [31:0] lo,
    output reg div0, 
);



endmodule;